module And(a,b,out);
input wire a,b;
output out;

assign out = a & b;

endmodule